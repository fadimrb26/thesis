* Define MOSFET models
.model PMOS PMOS (VTO=-0.4 KP=100u)
.model NMOS NMOS (VTO=0.4 KP=200u)
.model SWMODEL SW(Ron=1 Roff=1G Von=1 Voff=0.5)

* Power supply
Vdd VDD 0 1.1V

* Random noise source at input
Vnoise IN 0 PULSE(0 1u 0n 0.1n 0.1n 10n 30n)

* Inverter 1
M1 Q  N1 VDD VDD PMOS W=360n L=45n
M2 Q  N1 0   0   NMOS W=180n L=45n

* Inverter 2
M3 Qb N2 VDD VDD PMOS W=360n L=45n
M4 Qb N2 0   0   NMOS W=180n L=45n

* Capacitors at the outputs
C1 Q  0 100f  
C2 Qb 0 100f
C3 N1 0 100f
C4 N2 0 100f  

* Switch to connect input to the latch
S1 Qb IN CLK 0 SWMODEL
S2 Qb N1 CLK 0 SWMODEL
S3 Q  N2 CLK 0 SWMODEL
S4 Q  N1 NCLK 0 SWMODEL
S5 Qb N2 NCLK 0 SWMODEL  

* Clock signals (CLK high for 10ns, low for 20ns)
Vclk CLK 0 PULSE(0 1.8 0n 0.1n 0.1n 10n 30n)  
Vnclk NCLK 0 PULSE(1.8 0 0n 0.1n 0.1n 10n 30n) 

* Simulation control
.tran 0.1n 60n

.end
