* Define MOSFET models
.model PMOS PMOS (VTO=-0.4 KP=100u)
.model NMOS NMOS (VTO=0.4 KP=200u)
.model SWMODEL SW(Ron=1 Roff=1G Von=1 Voff=0.5)

* Define the latch subcircuit with initialization parameters
.SUBCKT LATCH Q Qb VDD GND PARAMS: VQ_init=0 VQb_init=0
* Inverter 1
M1 Q  Qb VDD VDD PMOS W=360n L=45n
M2 Q  Qb GND GND NMOS W=180n L=45n

* Inverter 2
M3 Qb Q VDD VDD PMOS W=360n L=45n
M4 Qb Q GND GND NMOS W=180n L=45n

* Capacitors at the outputs
C1 Q  GND 100f  
C2 Qb GND 100f

* Set initial conditions using parameters
.IC V(Q)={VQ_init} V(Qb)={VQb_init}
.ENDS LATCH

* Power supply
Vdd VDD 0 1.1V

* Instantiate the latches
X0 Q0 Qb0 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X1 Q4 Qb4 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X2 Q4 Qb4 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X3 Q4 Qb4 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X4 Q0 Qb0 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X5 Q3 Qb3 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X6 Q4 Qb4 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X7 Q0 Qb0 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X8 Q1 Qb1 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X9 Q4 Qb4 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X10 Q2 Qb2 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X11 Q2 Qb2 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0
X12 Q2 Qb2 VDD 0 LATCH PARAMS: VQ_init=0 VQb_init=0

* Connection between latch 0 and latches 1, 2, 3, and 4
* Latch 0 to Latch 1
S0_01 Q0 N0 FLY_CTRL0 0 SWMODEL
S1_01 Q1 N1 FLY_CTRL0 0 SWMODEL
S2_01 Qb0 N2 FLY_CTRL0 0 SWMODEL
S3_01 Qb1 N3 FLY_CTRL0 0 SWMODEL

S0i_01 Qb0 N0 NFLY_CTRL0 0 SWMODEL
S1i_01 Q1 N1 NFLY_CTRL0 0 SWMODEL
S2i_01 Q0 N2 NFLY_CTRL0 0 SWMODEL
S3i_01 Qb1 N3 NFLY_CTRL0 0 SWMODEL

* Latch 0 to Latch 2
S0_02 Q0 N4 FLY_CTRL1 0 SWMODEL
S1_02 Q2 N5 FLY_CTRL1 0 SWMODEL
S2_02 Qb0 N6 FLY_CTRL1 0 SWMODEL
S3_02 Qb2 N7 FLY_CTRL1 0 SWMODEL

S0i_02 Qb0 N4 NFLY_CTRL1 0 SWMODEL
S1i_02 Q2 N5 NFLY_CTRL1 0 SWMODEL
S2i_02 Q0 N6 NFLY_CTRL1 0 SWMODEL
S3i_02 Qb2 N7 NFLY_CTRL1 0 SWMODEL

* Latch 0 to Latch 3
S0_03 Q0 N8 FLY_CTRL2 0 SWMODEL
S1_03 Q3 N9 FLY_CTRL2 0 SWMODEL
S2_03 Qb0 N10 FLY_CTRL2 0 SWMODEL
S3_03 Qb3 N11 FLY_CTRL2 0 SWMODEL

S0i_03 Qb0 N8 NFLY_CTRL2 0 SWMODEL
S1i_03 Q3 N9 NFLY_CTRL2 0 SWMODEL
S2i_03 Q0 N10 NFLY_CTRL2 0 SWMODEL
S3i_03 Qb3 N11 NFLY_CTRL2 0 SWMODEL

* Latch 0 to Latch 4
S0_04 Q0 N12 FLY_CTRL3 0 SWMODEL
S1_04 Q4 N13 FLY_CTRL3 0 SWMODEL
S2_04 Qb0 N14 FLY_CTRL3 0 SWMODEL
S3_04 Qb4 N15 FLY_CTRL3 0 SWMODEL

S0i_04 Qb0 N12 NFLY_CTRL3 0 SWMODEL
S1i_04 Q4 N13 NFLY_CTRL3 0 SWMODEL
S2i_04 Q0 N14 NFLY_CTRL3 0 SWMODEL
S3i_04 Qb4 N15 NFLY_CTRL3 0 SWMODEL

* Connection between latch 1 and latches 2, 3, and 4
* Latch 1 to Latch 2
S0_12 Q1 N16 FLY_CTRL4 0 SWMODEL
S1_12 Q2 N17 FLY_CTRL4 0 SWMODEL
S2_12 Qb1 N18 FLY_CTRL4 0 SWMODEL
S3_12 Qb2 N19 FLY_CTRL4 0 SWMODEL

S0i_12 Qb1 N16 NFLY_CTRL4 0 SWMODEL
S1i_12 Q2 N17 NFLY_CTRL4 0 SWMODEL
S2i_12 Q1 N18 NFLY_CTRL4 0 SWMODEL
S3i_12 Qb2 N19 NFLY_CTRL4 0 SWMODEL

* Latch 1 to Latch 3
S0_13 Q1 N20 FLY_CTRL5 0 SWMODEL
S1_13 Q3 N21 FLY_CTRL5 0 SWMODEL
S2_13 Qb1 N22 FLY_CTRL5 0 SWMODEL
S3_13 Qb3 N23 FLY_CTRL5 0 SWMODEL

S0i_13 Qb1 N20 NFLY_CTRL5 0 SWMODEL
S1i_13 Q3 N21 NFLY_CTRL5 0 SWMODEL
S2i_13 Q1 N22 NFLY_CTRL5 0 SWMODEL
S3i_13 Qb3 N23 NFLY_CTRL5 0 SWMODEL

* Latch 1 to Latch 4
S0_14 Q1 N24 FLY_CTRL6 0 SWMODEL
S1_14 Q4 N25 FLY_CTRL6 0 SWMODEL
S2_14 Qb1 N26 FLY_CTRL6 0 SWMODEL
S3_14 Qb4 N27 FLY_CTRL6 0 SWMODEL

S0i_14 Qb1 N24 NFLY_CTRL6 0 SWMODEL
S1i_14 Q4 N25 NFLY_CTRL6 0 SWMODEL
S2i_14 Q1 N26 NFLY_CTRL6 0 SWMODEL
S3i_14 Qb4 N27 NFLY_CTRL6 0 SWMODEL

* Latch 2 to Latch 4
S0_24 Q2 N32 FLY_CTRL8 0 SWMODEL
S1_24 Q4 N33 FLY_CTRL8 0 SWMODEL
S2_24 Qb2 N34 FLY_CTRL8 0 SWMODEL
S3_24 Qb4 N35 FLY_CTRL8 0 SWMODEL

S0i_24 Qb2 N32 NFLY_CTRL8 0 SWMODEL
S1i_24 Q4 N33 NFLY_CTRL8 0 SWMODEL
S2i_24 Q2 N34 NFLY_CTRL8 0 SWMODEL
S3i_24 Qb4 N35 NFLY_CTRL8 0 SWMODEL
* Flying capacitors
C_fly_0 N0 N1 20f
C_fly_1 N2 N3 20f
C_fly_2 N4 N5 20f
C_fly_3 N6 N7 20f

C_fly_4 N8 N9 20f
C_fly_5 N10 N11 20f

C_fly_6 N12 N13 20f
C_fly_7 N14 N15 20f

C_fly_8 N16 N17 20f
C_fly_9 N18 N19 20f

C_fly_10 N20 N21 20f
C_fly_11 N22 N23 20f

C_fly_12 N24 N25 20f
C_fly_13 N26 N27 20f 

C_fly_14 N28 N29 20f
C_fly_15 N30 N31 20f

C_fly_16 N32 N33 20f
C_fly_17 N34 N35 20f
* Control signals for flying capacitors
Vfly_ctrl0 FLY_CTRL0 0 DC 0
Vnfly_ctrl0 NFLY_CTRL0 0 DC 1.1

Vfly_ctrl1 FLY_CTRL1 0 DC 0
Vnfly_ctrl1 NFLY_CTRL1 0 DC 1.1

Vfly_ctrl2 FLY_CTRL2 0 DC 0
Vnfly_ctrl2 NFLY_CTRL2 0 DC 1.1

Vfly_ctrl3 FLY_CTRL3 0 DC 0
Vnfly_ctrl3 NFLY_CTRL3 0 DC 1.1

Vfly_ctrl4 FLY_CTRL4 0 DC 0
Vnfly_ctrl4 NFLY_CTRL4 0 DC 1.1

Vfly_ctrl5 FLY_CTRL5 0 DC 0
Vnfly_ctrl5 NFLY_CTRL5 0 DC 1.1

Vfly_ctrl6 FLY_CTRL6 0 DC 0
Vnfly_ctrl6 NFLY_CTRL6 0 DC 1.1

Vfly_ctrl7 FLY_CTRL7 0 DC 0
Vnfly_ctrl7 NFLY_CTRL7 0 DC 1.1

Vfly_ctrl8 FLY_CTRL8 0 DC 0
Vnfly_ctrl8 NFLY_CTRL8 0 DC 1.1
* Simulation control
.tran 0.1n 120n

.end
